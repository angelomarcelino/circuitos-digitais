library verilog;
use verilog.vl_types.all;
entity Counter2_VHDL_vlg_vec_tst is
end Counter2_VHDL_vlg_vec_tst;
