library verilog;
use verilog.vl_types.all;
entity demux_vlg_vec_tst is
end demux_vlg_vec_tst;
