library verilog;
use verilog.vl_types.all;
entity Counter2_VHDL_vlg_check_tst is
    port(
        Output          : in     vl_logic_vector(0 to 6);
        sampler_rx      : in     vl_logic
    );
end Counter2_VHDL_vlg_check_tst;
